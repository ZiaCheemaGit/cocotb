-- Copyright cocotb contributors
-- Licensed under the Revised BSD License, see LICENSE for details.
-- SPDX-License-Identifier: BSD-3-Clause

library ieee;
use ieee.std_logic_1164.all;

entity vhdl_top_a is
end vhdl_top_a;

architecture rtl of vhdl_top_a is
    signal flag : std_logic := '0';
begin
end rtl;

entity vhdl_top_b is
end vhdl_top_b;

architecture rtl of vhdl_top_b is
    signal flag : std_logic := '0';
begin
end rtl;
