// Copyright cocotb contributors
// Licensed under the Revised BSD License, see LICENSE for details.
// SPDX-License-Identifier: BSD-3-Clause

module verilog_top_a;
    reg flag = 0;
endmodule

module verilog_top_b;
    reg flag = 0;
endmodule
